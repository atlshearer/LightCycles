PACKAGE Game IS
  TYPE t_LocationState IS (Empty, Player1, Player2, Path);
END PACKAGE;